`timescale 1ns/1ps

module alu(opcode, inA, inB,in_apsr, out, out_apsr, branch_con);

input [3:0] opcode;
input [15:0] inA, inB, in_apsr;
output reg [15:0] out, out_apsr;
output reg branch_con; 

localparam  push=0, pop=1, sub_sp=2, cmp=3, movs=4, mov=5, ldr=6, str=7, 
            ldr_nop=8, add_sp=9, branch_nc= 10, adds_3op=11, branch_c=12, strb=13, ldrb=14, adds_2op=15;

`define in_carry in_apsr[1]
`define in_zero in_apsr[2]
`define in_overflow in_apsr[0]
`define in_negative in_apsr[3]


`define out_overflow out_apsr[0]
`define out_carry out_apsr[1]
`define out_zero out_apsr[2]
`define out_negative out_apsr[3]

always @(opcode, inA, inB) begin
	branch_con = 1'b0;
	case(opcode)
	push: begin //inA= Stack Pointer  
		out <= inA-1;
		`out_carry = `in_carry ;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_zero = `in_zero ; 
		$display("PUSH");
	      end 

	pop: begin
		//SP increment 
		
		//SP increase by 2 as registers both are being poped
		$display("POP");
	     end

	sub_sp: begin
//		 out = inA - inB;
		 //if(out==0) `out_zero = 0;
		 out = inA - inB ; 
		if(out==0) `out_zero = 1'b1 ;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_carry = `in_carry ;
		$display("ALU SUB inA: %h  inB: %h out:%h", inA, inB, out);
	     end
	
	add_sp: begin
		{`out_overflow, out} = inA + inB; 
		$display("ALU ADD inA: %h  inB: %h out:%h", inA, inB, out);
	     end
   
        adds_2op: begin
		{`out_overflow, out} = inA + inB + `in_carry; 
		$display("ALU ADD 2OP inA: %h  inB: %h out:%h", inA, inB, out);
	     end
      
        adds_3op: begin
		{`out_overflow, out} = inA + inB; 
		$display("ALU ADD inA: %h  inB: %h out:%h", inA, inB, out);
	     end
       
	cmp: begin
		 out= inA-inB;
		 if(out==0) `out_zero = 1'b1 ;
		 else `out_zero = 1'b0 ;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_carry = `in_carry ;
		$display("CMP inA=%h inB=%h ZF=%b",inA, inB, `out_zero);
	     end
	
	str: begin
	     end

	ldr: begin
	     end

	branch_c: begin
		if(`in_zero) begin
			out=inA;
			`out_zero= 1'b0;
			branch_con = 1'b1;
		end
                else `out_zero= `in_zero;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_carry = `in_carry ;
	     end

	branch_nc: begin
		out=inA;
		
	    end

	movs: begin
		out= inA + inB;
		`out_carry = `in_carry ;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_zero = `in_zero ;
		$display("ALU MOVS inA: %h  inB: %h out:%h", inA, inB, out);
	     end

	mov: begin
		out= inB;
		`out_carry = `in_carry ;
		`out_overflow = `in_overflow ;
		`out_negative = `in_negative ;
		`out_zero = `in_zero ;
		$display("ALU MOV inA: %h  inB: %h out:%h", inA, inB, out);
	end


	endcase

end 

endmodule

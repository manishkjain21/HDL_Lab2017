`timescale 10ns/1ns

module cpu();

reg [15:0]addr;





endmodule

